module ver;
   initial $display("I am version 1");
endmodule
