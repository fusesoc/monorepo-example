module top;
   ver ver();
endmodule
