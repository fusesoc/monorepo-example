module ver;
   initial $display("I am version 2");
endmodule
